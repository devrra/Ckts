*** SPICE deck for cell simpleCS{sch} from library Common_Source
*** Created on Sat Aug 01, 2020 06:32:17
*** Last revised on Sat Aug 01, 2020 15:48:03
*** Written on Sat Aug 01, 2020 15:48:08 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: simpleCS{sch}
Mnmos@0 out b gnd gnd NMOS L=0.13U W=0.13U

* Spice Code nodes in cell cell 'simpleCS{sch}'
.include C:\Users\Yash Raj\Documents\electric\130nm.cir
Rd vdd out 16k
R1 vdd b 100k
R2 b 0 200k
Cin in b 0.1uF
Vvdd vdd 0 1.2
Vin in 0 sin(0 50m 10k)
.tran 10u 0.5m
.END
