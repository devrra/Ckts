*** SPICE deck for cell degeneratedCG{sch} from library CommonGate
*** Created on Tue Aug 04, 2020 15:24:42
*** Last revised on Tue Aug 04, 2020 16:40:52
*** Written on Tue Aug 04, 2020 16:40:58 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: degeneratedCG{sch}
Mnmos@0 out b s gnd NMOS L=0.13U W=0.13U

* Spice Code nodes in cell cell 'degeneratedCG{sch}'
.include C:\Users\Yash Raj\Documents\electric\130nm.cir
Vvdd vdd 0 1.2
Rs s a 10k
R1 vdd b 100k
R2 b 0 100k
R3 vdd a 300k
R4 a 0 100k
Cin in a 0.1uF
Vin in 0 sin(0 50m 10k)
.tran 10u .5m
.END
